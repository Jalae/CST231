///////////////////////////////////////////////////////////////////////////////
//Kehnin Dyer
//20120208
//Homework 2
//
///////////////////////////////////////////////////////////////////////////////
module Adder
(
	input		[5:0]	A,
						B,
	output	reg	[5:0]	C//,
//	output	reg		O
);
wire cout;
always@(*)
begin
C = A[5:0] + B[5:0];
//O = ((A[5]&B[5])|(~A[5]&~B[5]))^C[5];
end

endmodule

