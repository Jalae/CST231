
module Elevator_ButtonDecode(
	input	
	
);



endmodule

