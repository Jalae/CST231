

module SetDestination(

);


endmodule

